module vsync(
	input line_clk, 
	output vsync_out, 
	output blank_out
	);
   
   reg [10:0] count = 10'b0000000000;
   reg vsync  = 0;
   reg blank  = 0;

   always @(posedge line_clk)
	 if (count < 666)
	   count <= count + 1;
	 else
	   count <= 0;
   
   always @(posedge line_clk)
	 if (count < 600)
	   blank 		<= 0;
	 else
	   blank 		<= 1;
      
   always @(posedge line_clk)
	 begin
		if (count < 637)
		  vsync 	<= 1;
		else if (count >= 637 && count < 643)
		  vsync 	<= 0;
		else if (count >= 643)
		  vsync 	<= 1;
	 end

   assign vsync_out  = vsync;
   assign blank_out  = blank;
   
endmodule // hsync   

module hsync(
	input clk50, 
	output hsync_out, 
	output blank_out, 
	output newline_out
	);
   
   reg [10:0] count = 10'b0000000000;
   reg hsync 	= 0;
   reg blank 	= 0;
   reg newline 	= 0;

   always @(posedge clk50)
	 begin
		if (count < 1040)
		  count  <= count + 1;
		else
		  count  <= 0;
	 end
   
   always @(posedge clk50)
	 begin
		if (count == 0)
		  newline <= 1;
		else
		  newline <= 0;
	 end

   always @(posedge clk50)
	 begin
		if (count >= 800)
		  blank  <= 1;
		else
		  blank  <= 0;
	 end

   always @(posedge clk50)
	 begin
		if (count < 856) // pixel data plus front porch
		  hsync <= 1;
		else if (count >= 856 && count < 976)
		  hsync <= 0;
		else if (count >= 976)
		  hsync <= 1;
	 end // always @ (posedge clk50)
				 
   assign hsync_out    = hsync;
   assign blank_out    = blank;
   assign newline_out  = newline;
   
endmodule // hsync


module color(
	input clk, 
	input blank, 
	output [7:0] red_out, 
	output [7:0] green_out, 
	output [7:0] blue_out
	);
	
   reg [8:0] count;
   
   always @(posedge clk)
	 begin
		if (blank)
		  count 	<= 0;
		else
		  count 	<= 1;
	 end

   assign red_out	 = (blank) ? 0 : 8'b11111111;
	assign green_out = (blank) ? 0 : 8'b01111111;
	assign blue_out  = (blank) ? 0 : 8'b00001111;
   
endmodule // color

module gridandwave(
	input clk, 
	input blank, 
	input hsync,
	input vsync,
	input cursorX_EN,
	input cursorY_EN,
	input [10:0] cursorY1,
	input [10:0] cursorY2,
	input [10:0] cursorX1,
	input [10:0] cursorX2,
	input [13:0] waveSigIn1,
	input [13:0] waveSigIn2,
	input [10:0] wave1YOffset,
	input [10:0] wave2YOffset,	
	input waveSigIn1_En,
	input waveSigIn2_En,
	output [7:0] red_out, 
	output [7:0] green_out, 
	output [7:0] blue_out,
	output [10:0] sX,
	output [10:0] sY
	);
	localparam gridoffset = 20;
	reg [19:0] x;
	reg [19:0] y;
   reg [8:0] count;
   reg [7:0] pixel_R = 0;
	reg [7:0] pixel_G = 0;
	reg [7:0] pixel_B = 0;
	reg [8:0] i;
	assign sX = x;
	assign sY = y;
   always @(posedge clk)
	 begin
		if (blank) begin
			if(hsync) begin
			x <= 0;
			end else if (vsync) begin
			x <= 0;
			end
		end else begin
			x <= x+1;
			//wave code
			if (waveSigIn1_En && y == (waveSigIn1 + wave1YOffset)) begin
			pixel_R <= 8'b00000000;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if (waveSigIn2_En && (y == waveSigIn2 + wave2YOffset)) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b00000000;
			pixel_B <= 8'b11111111;
			//cursor code
			end else if(cursorX_EN && x == cursorX1) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b00000000;
			end else if (cursorX_EN && x == cursorX2) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b00000000;
			end else if (cursorY_EN && y == cursorY1) begin
			pixel_R <= 8'b00000000;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b00000000;
			end else if (cursorY_EN && y == cursorY2) begin
			pixel_R <= 8'b00000000;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b00000000;
			//grid
			end else if(y == 60 * 1) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(y == 60 * 2) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(y == 60 * 3) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(y == 60 * 4) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(y == 60 * 5) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(y == 60 * 6) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(y == 60 * 7) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(y == 60 * 8) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(y == 60 * 9) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			//X Grid
			end else if(x == (60 * 1) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 2) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 3) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 4) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 5) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 6) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 7) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 8) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 9) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 10) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 11) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 12) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 13) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else if(x == (60 * 14) - gridoffset) begin
			pixel_R <= 8'b11111111;
			pixel_G <= 8'b11111111;
			pixel_B <= 8'b11111111;
			end else begin
			pixel_R <= 8'b0;
			pixel_G <= 8'b0;
			pixel_B <= 8'b0;
			end
		end
	 end
	
	always @(posedge hsync) begin
		if(vsync) begin
			y <= 0;
		end else begin
			y <= y + 1;
		end
	end
   assign red_out	 = (blank) ? 0 : pixel_R;
	assign green_out = (blank) ? 0 : pixel_G;
	assign blue_out  = (blank) ? 0 : pixel_B;
   
endmodule // color