/* Top level modile for FPGA_MiniProject
Alexander Bolton - 200938078
Haider Shafiq - 201207577
N-Channel Oscilloscope */

module FPGA_MiniProject





endmodule 