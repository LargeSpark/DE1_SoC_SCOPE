/* Measurements for Scope
 * DE1-SoC Scope, FPGA Mini-Project
 *	Alexander Bolton & Haider Shafiq
 */
 
 module Scope_Measurements 
 (
 
 
 )