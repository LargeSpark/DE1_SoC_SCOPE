module Measure(
	input  c1x,
	input  c2x,
	input  c1y,
	input  c2y,
	output xD,
	output yD
);
// Register to store initial number i.e. = 500mV
reg [5:0] num = 0;


endmodule 